library verilog;
use verilog.vl_types.all;
entity alsu_tb is
end alsu_tb;
